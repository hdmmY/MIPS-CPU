`timescale 1ns / 1ps
/**
 * @module ins_mem.v
 * @brief instruction cache memory (ROM)
 * @param DATA_WIDTH data width
 * @param BUS_WIDTH bus width
 * @param CODE_FILE MIPS assembly hexdecimal code file
 * @input addr memory address
 * @output rdata instruction read out from memory
 */
 module ins_mem
 #(parameter DATA_WIDTH = 32, BUS_WIDTH = 10, CODE_FILE= "D:/benchmark.hex")
 (
 	input [BUS_WIDTH-1:0] addr,
 	output [DATA_WIDTH-1:0] rdata
 );

 	reg [DATA_WIDTH-1:0] ROM [0:(2**BUS_WIDTH)-1];

 	initial begin
 	ROM[0] = 32'h20110001;
     ROM[1] = 32'h08000c05;
     ROM[2] = 32'h20110001;
     ROM[3] = 32'h20120002;
     ROM[4] = 32'h20130003;
     ROM[5] = 32'h08000c09;
     ROM[6] = 32'h20110001;
     ROM[7] = 32'h20120002;
     ROM[8] = 32'h20130003;
     ROM[9] = 32'h08000c0d;
     ROM[10] = 32'h20110001;
     ROM[11] = 32'h20120002;
     ROM[12] = 32'h20130003;
     ROM[13] = 32'h08000c11;
     ROM[14] = 32'h20110001;
     ROM[15] = 32'h20120002;
     ROM[16] = 32'h20130003;
     ROM[17] = 32'h0c000cb8;
     ROM[18] = 32'h20100001;
     ROM[19] = 32'h20110001;
     ROM[20] = 32'h00118fc0;
     ROM[21] = 32'h00112020;
     ROM[22] = 32'h20020022;
     ROM[23] = 32'h0000000c;
     ROM[24] = 32'h00118882;
     ROM[25] = 32'h12200001;
     ROM[26] = 32'h08000c15;
     ROM[27] = 32'h00112020;
     ROM[28] = 32'h20020022;
     ROM[29] = 32'h0000000c;
     ROM[30] = 32'h20110001;
     ROM[31] = 32'h00118880;
     ROM[32] = 32'h00112020;
     ROM[33] = 32'h20020022;
     ROM[34] = 32'h0000000c;
     ROM[35] = 32'h12200001;
     ROM[36] = 32'h08000c1f;
     ROM[37] = 32'h20110001;
     ROM[38] = 32'h00118fc0;
     ROM[39] = 32'h00112020;
     ROM[40] = 32'h20020022;
     ROM[41] = 32'h0000000c;
     ROM[42] = 32'h001188c3;
     ROM[43] = 32'h00112020;
     ROM[44] = 32'h20020022;
     ROM[45] = 32'h0000000c;
     ROM[46] = 32'h00118903;
     ROM[47] = 32'h00112020;
     ROM[48] = 32'h20020022;
     ROM[49] = 32'h0000000c;
     ROM[50] = 32'h00118903;
     ROM[51] = 32'h00112020;
     ROM[52] = 32'h20020022;
     ROM[53] = 32'h0000000c;
     ROM[54] = 32'h00118903;
     ROM[55] = 32'h00112020;
     ROM[56] = 32'h20020022;
     ROM[57] = 32'h0000000c;
     ROM[58] = 32'h00118903;
     ROM[59] = 32'h00112020;
     ROM[60] = 32'h20020022;
     ROM[61] = 32'h0000000c;
     ROM[62] = 32'h00118903;
     ROM[63] = 32'h00112020;
     ROM[64] = 32'h20020022;
     ROM[65] = 32'h0000000c;
     ROM[66] = 32'h00118903;
     ROM[67] = 32'h00112020;
     ROM[68] = 32'h20020022;
     ROM[69] = 32'h0000000c;
     ROM[70] = 32'h00118903;
     ROM[71] = 32'h00112020;
     ROM[72] = 32'h20020022;
     ROM[73] = 32'h0000000c;
     ROM[74] = 32'h20100001;
     ROM[75] = 32'h00109fc0;
     ROM[76] = 32'h00139fc3;
     ROM[77] = 32'h00008021;
     ROM[78] = 32'h2012000c;
     ROM[79] = 32'h24160003;
     ROM[80] = 32'h26100001;
     ROM[81] = 32'h3210000f;
     ROM[82] = 32'h20080008;
     ROM[83] = 32'h20090001;
     ROM[84] = 32'h00139900;
     ROM[85] = 32'h02709825;
     ROM[86] = 32'h00132020;
     ROM[87] = 32'h20020022;
     ROM[88] = 32'h0000000c;
     ROM[89] = 32'h01094022;
     ROM[90] = 32'h1500fff9;
     ROM[91] = 32'h22100001;
     ROM[92] = 32'h2018000f;
     ROM[93] = 32'h02188024;
     ROM[94] = 32'h00108700;
     ROM[95] = 32'h20080008;
     ROM[96] = 32'h20090001;
     ROM[97] = 32'h00139902;
     ROM[98] = 32'h02709825;
     ROM[99] = 32'h00132021;
     ROM[100] = 32'h20020022;
     ROM[101] = 32'h0000000c;
     ROM[102] = 32'h01094022;
     ROM[103] = 32'h1500fff9;
     ROM[104] = 32'h00108702;
     ROM[105] = 32'h02c9b022;
     ROM[106] = 32'h12c00001;
     ROM[107] = 32'h08000c50;
     ROM[108] = 32'h00004020;
     ROM[109] = 32'h01084027;
     ROM[110] = 32'h00084400;
     ROM[111] = 32'h3508ffff;
     ROM[112] = 32'h00082021;
     ROM[113] = 32'h20020022;
     ROM[114] = 32'h0000000c;
     ROM[115] = 32'h2010ffff;
     ROM[116] = 32'h20110000;
     ROM[117] = 32'hae300000;
     ROM[118] = 32'h22100001;
     ROM[119] = 32'h22310004;
     ROM[120] = 32'hae300000;
     ROM[121] = 32'h22100001;
     ROM[122] = 32'h22310004;
     ROM[123] = 32'hae300000;
     ROM[124] = 32'h22100001;
     ROM[125] = 32'h22310004;
     ROM[126] = 32'hae300000;
     ROM[127] = 32'h22100001;
     ROM[128] = 32'h22310004;
     ROM[129] = 32'hae300000;
     ROM[130] = 32'h22100001;
     ROM[131] = 32'h22310004;
     ROM[132] = 32'hae300000;
     ROM[133] = 32'h22100001;
     ROM[134] = 32'h22310004;
     ROM[135] = 32'hae300000;
     ROM[136] = 32'h22100001;
     ROM[137] = 32'h22310004;
     ROM[138] = 32'hae300000;
     ROM[139] = 32'h22100001;
     ROM[140] = 32'h22310004;
     ROM[141] = 32'hae300000;
     ROM[142] = 32'h22100001;
     ROM[143] = 32'h22310004;
     ROM[144] = 32'hae300000;
     ROM[145] = 32'h22100001;
     ROM[146] = 32'h22310004;
     ROM[147] = 32'hae300000;
     ROM[148] = 32'h22100001;
     ROM[149] = 32'h22310004;
     ROM[150] = 32'hae300000;
     ROM[151] = 32'h22100001;
     ROM[152] = 32'h22310004;
     ROM[153] = 32'hae300000;
     ROM[154] = 32'h22100001;
     ROM[155] = 32'h22310004;
     ROM[156] = 32'hae300000;
     ROM[157] = 32'h22100001;
     ROM[158] = 32'h22310004;
     ROM[159] = 32'hae300000;
     ROM[160] = 32'h22100001;
     ROM[161] = 32'h22310004;
     ROM[162] = 32'hae300000;
     ROM[163] = 32'h22100001;
     ROM[164] = 32'h22310004;
     ROM[165] = 32'h22100001;
     ROM[166] = 32'h00008020;
     ROM[167] = 32'h2011003c;
     ROM[168] = 32'h8e130000;
     ROM[169] = 32'h8e340000;
     ROM[170] = 32'h0274402a;
     ROM[171] = 32'h11000002;
     ROM[172] = 32'hae330000;
     ROM[173] = 32'hae140000;
     ROM[174] = 32'h2231fffc;
     ROM[175] = 32'h1611fff8;
     ROM[176] = 32'h00102020;
     ROM[177] = 32'h20020022;
     ROM[178] = 32'h0000000c;
     ROM[179] = 32'h22100004;
     ROM[180] = 32'h2011003c;
     ROM[181] = 32'h1611fff2;
     ROM[182] = 32'h2002000a;
     ROM[183] = 32'h0000000c;
     ROM[184] = 32'h20100000;
     ROM[185] = 32'h22100001;
     ROM[186] = 32'h00102020;
     ROM[187] = 32'h20020022;
     ROM[188] = 32'h0000000c;
     ROM[189] = 32'h22100002;
     ROM[190] = 32'h00102020;
     ROM[191] = 32'h20020022;
     ROM[192] = 32'h0000000c;
     ROM[193] = 32'h22100003;
     ROM[194] = 32'h00102020;
     ROM[195] = 32'h20020022;
     ROM[196] = 32'h0000000c;
     ROM[197] = 32'h22100004;
     ROM[198] = 32'h00102020;
     ROM[199] = 32'h20020022;
     ROM[200] = 32'h0000000c;
     ROM[201] = 32'h22100005;
     ROM[202] = 32'h00102020;
     ROM[203] = 32'h20020022;
     ROM[204] = 32'h0000000c;
     ROM[205] = 32'h22100006;
     ROM[206] = 32'h00102020;
     ROM[207] = 32'h20020022;
     ROM[208] = 32'h0000000c;
     ROM[209] = 32'h22100007;
     ROM[210] = 32'h00102020;
     ROM[211] = 32'h20020022;
     ROM[212] = 32'h0000000c;
     ROM[213] = 32'h22100008;
     ROM[214] = 32'h00102020;
     ROM[215] = 32'h20020022;
     ROM[216] = 32'h20020022;
     ROM[217] = 32'h0000000c;
     ROM[218] = 32'h03e00008;
 	end
 	assign rdata = ROM[addr];
 endmodule