module hellow_world;

initial begin
    $display("Hello World by hdm.");
    #10 $finish;
end

endmodule // hellow_world